/*******************************************************************************
Creator:        Hai Cao Xuan (caoxuanhaipr@gmail.com)

Additional Contributions by:

File Name:      my_pkg.svh
Design Name:    My Package
Project Name:   Computer Architecture Examples
Description:    Package of configuration and defines

Changelog:      06.07.2022 - First draft, v0.1

********************************************************************************
Copyright (c) 2022 Hai Cao Xuan
*******************************************************************************/

package my_pkg;


endpackage : my_pkg
